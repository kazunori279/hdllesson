/*

  rom.v
  
  Represents an instruction rom for debug purpose.
  
  */

`include "src/defines.v"

module rom (
	input [`WORD] pc,
	output reg [`WORD] inst
);

	always_comb begin
		case (pc)
		
32'd0: inst = 32'h00000000;
32'd4: inst = 32'h00000000;
32'd8: inst = 32'h00000000;
32'd12: inst = 32'h00000000;
32'd16: inst = 32'h00000000;
32'd20: inst = 32'h00000000;
32'd24: inst = 32'h00000000;
32'd28: inst = 32'h00000000;
32'd32: inst = 32'h00000000;
32'd36: inst = 32'h00000000;
32'd40: inst = 32'h00000000;
32'd44: inst = 32'h2008ffff;
32'd48: inst = 32'hac080000;
32'd52: inst = 32'h20080001;
32'd56: inst = 32'ha4080000;
32'd60: inst = 32'h8c090000;
32'd64: inst = 32'h3c0fffff;
32'd68: inst = 32'h35ef0001;
32'd72: inst = 32'h152ffffc;
32'd76: inst = 32'h00000000;
32'd80: inst = 32'h00000000;
32'd84: inst = 32'h2008ffff;
32'd88: inst = 32'hac080000;
32'd92: inst = 32'h20080001;
32'd96: inst = 32'ha4080002;
32'd100: inst = 32'h8c090000;
32'd104: inst = 32'h3c0f0001;
32'd108: inst = 32'h35efffff;
32'd112: inst = 32'h152ffffc;
32'd116: inst = 32'h00000000;
32'd120: inst = 32'h00000000;
32'd124: inst = 32'h2008ffff;
32'd128: inst = 32'hac080000;
32'd132: inst = 32'h20080001;
32'd136: inst = 32'ha0080000;
32'd140: inst = 32'h8c090000;
32'd144: inst = 32'h3c0fffff;
32'd148: inst = 32'h35efff01;
32'd152: inst = 32'h152ffffc;
32'd156: inst = 32'h00000000;
32'd160: inst = 32'h00000000;
32'd164: inst = 32'h2008ffff;
32'd168: inst = 32'hac080000;
32'd172: inst = 32'h20080001;
32'd176: inst = 32'ha0080001;
32'd180: inst = 32'h8c090000;
32'd184: inst = 32'h3c0fffff;
32'd188: inst = 32'h35ef01ff;
32'd192: inst = 32'h152ffffc;
32'd196: inst = 32'h00000000;
32'd200: inst = 32'h00000000;
32'd204: inst = 32'h2008ffff;
32'd208: inst = 32'hac080000;
32'd212: inst = 32'h20080001;
32'd216: inst = 32'ha0080002;
32'd220: inst = 32'h8c090000;
32'd224: inst = 32'h3c0fff01;
32'd228: inst = 32'h35efffff;
32'd232: inst = 32'h152ffffc;
32'd236: inst = 32'h00000000;
32'd240: inst = 32'h00000000;
32'd244: inst = 32'h2008ffff;
32'd248: inst = 32'hac080000;
32'd252: inst = 32'h20080001;
32'd256: inst = 32'ha0080003;
32'd260: inst = 32'h8c090000;
32'd264: inst = 32'h3c0f01ff;
32'd268: inst = 32'h35efffff;
32'd272: inst = 32'h152ffffc;
32'd276: inst = 32'h00000000;
32'd280: inst = 32'h00000000;
32'd284: inst = 32'h3c080102;
32'd288: inst = 32'h3508f3f4;
32'd292: inst = 32'hac080000;
32'd296: inst = 32'h94080000;
32'd300: inst = 32'h94090002;
32'd304: inst = 32'h200f0000;
32'd308: inst = 32'h35eff3f4;
32'd312: inst = 32'h150ffffd;
32'd316: inst = 32'h00000000;
32'd320: inst = 32'h200f0102;
32'd324: inst = 32'h152ffffe;
32'd328: inst = 32'h00000000;
32'd332: inst = 32'h00000000;
32'd336: inst = 32'h3c080102;
32'd340: inst = 32'h3508f3f4;
32'd344: inst = 32'hac080000;
32'd348: inst = 32'h84080000;
32'd352: inst = 32'h84090002;
32'd356: inst = 32'h200ff3f4;
32'd360: inst = 32'h150ffffe;
32'd364: inst = 32'h00000000;
32'd368: inst = 32'h200f0102;
32'd372: inst = 32'h152ffffe;
32'd376: inst = 32'h00000000;
32'd380: inst = 32'h00000000;
32'd384: inst = 32'h3c08f102;
32'd388: inst = 32'h3508f304;
32'd392: inst = 32'hac080000;
32'd396: inst = 32'h90080000;
32'd400: inst = 32'h90090001;
32'd404: inst = 32'h900a0002;
32'd408: inst = 32'h900b0003;
32'd412: inst = 32'h200f0004;
32'd416: inst = 32'h150ffffe;
32'd420: inst = 32'h00000000;
32'd424: inst = 32'h200f00f3;
32'd428: inst = 32'h152ffffe;
32'd432: inst = 32'h00000000;
32'd436: inst = 32'h200f0002;
32'd440: inst = 32'h154ffffe;
32'd444: inst = 32'h00000000;
32'd448: inst = 32'h200f00f1;
32'd452: inst = 32'h156ffffe;
32'd456: inst = 32'h00000000;
32'd460: inst = 32'h00000000;
32'd464: inst = 32'h3c08f102;
32'd468: inst = 32'h3508f304;
32'd472: inst = 32'hac080000;
32'd476: inst = 32'h80080000;
32'd480: inst = 32'h80090001;
32'd484: inst = 32'h800a0002;
32'd488: inst = 32'h800b0003;
32'd492: inst = 32'h200f0004;
32'd496: inst = 32'h150ffffe;
32'd500: inst = 32'h00000000;
32'd504: inst = 32'h200ffff3;
32'd508: inst = 32'h152ffffe;
32'd512: inst = 32'h00000000;
32'd516: inst = 32'h200f0002;
32'd520: inst = 32'h154ffffe;
32'd524: inst = 32'h00000000;
32'd528: inst = 32'h200ffff1;
32'd532: inst = 32'h156ffffe;
32'd536: inst = 32'h00000000;
32'd540: inst = 32'h00000000;
32'd544: inst = 32'h20080001;
32'd548: inst = 32'hac080000;
32'd552: inst = 32'h8c090000;
32'd556: inst = 32'h21ef0001;
32'd560: inst = 32'h152ffffe;
32'd564: inst = 32'h00000000;
32'd568: inst = 32'h00000000;
32'd572: inst = 32'h3c080001;
32'd576: inst = 32'h200f0001;
32'd580: inst = 32'h000f7c00;
32'd584: inst = 32'h150ffffd;
32'd588: inst = 32'h00000000;
32'd592: inst = 32'h00000000;
32'd596: inst = 32'h20080001;
32'd600: inst = 32'h3109ffff;
32'd604: inst = 32'h350affff;
32'd608: inst = 32'h390bffff;
32'd612: inst = 32'h200f0001;
32'd616: inst = 32'h152ffffe;
32'd620: inst = 32'h00000000;
32'd624: inst = 32'h3c0fffff;
32'd628: inst = 32'h000f7c02;
32'd632: inst = 32'h154ffffa;
32'd636: inst = 32'h00000000;
32'd640: inst = 32'h3c0ffffe;
32'd644: inst = 32'h000f7c02;
32'd648: inst = 32'h156ffff6;
32'd652: inst = 32'h00000000;
32'd656: inst = 32'h00000000;
32'd660: inst = 32'h20080001;
32'd664: inst = 32'h2909ffff;
32'd668: inst = 32'h2d0a0000;
32'd672: inst = 32'h1520ffff;
32'd676: inst = 32'h00000000;
32'd680: inst = 32'h1540fffd;
32'd684: inst = 32'h00000000;
32'd688: inst = 32'h00000000;
32'd692: inst = 32'h20080001;
32'd696: inst = 32'h21090001;
32'd700: inst = 32'h200f0002;
32'd704: inst = 32'h152ffffe;
32'd708: inst = 32'h00000000;
32'd712: inst = 32'h00000000;
32'd716: inst = 32'h24080001;
32'd720: inst = 32'h25090001;
32'd724: inst = 32'h200f0002;
32'd728: inst = 32'h152ffffe;
32'd732: inst = 32'h00000000;
32'd736: inst = 32'h00000000;
32'd740: inst = 32'h2008ffff;
32'd744: inst = 32'h19000003;
32'd748: inst = 32'h00000000;
32'd752: inst = 32'h080000ba;
32'd756: inst = 32'h00000000;
32'd760: inst = 32'h00000000;
32'd764: inst = 32'h20080001;
32'd768: inst = 32'h1d000003;
32'd772: inst = 32'h00000000;
32'd776: inst = 32'h080000c0;
32'd780: inst = 32'h00000000;
32'd784: inst = 32'h00000000;
32'd788: inst = 32'h2008ffff;
32'd792: inst = 32'h05000003;
32'd796: inst = 32'h00000000;
32'd800: inst = 32'h080000c6;
32'd804: inst = 32'h00000000;
32'd808: inst = 32'h00000000;
32'd812: inst = 32'h20080000;
32'd816: inst = 32'h05010003;
32'd820: inst = 32'h00000000;
32'd824: inst = 32'h080000cc;
32'd828: inst = 32'h00000000;
32'd832: inst = 32'h00000000;
32'd836: inst = 32'h04010003;
32'd840: inst = 32'h00000000;
32'd844: inst = 32'h080000d1;
32'd848: inst = 32'h00000000;
32'd852: inst = 32'h00000000;
32'd856: inst = 32'h10000003;
32'd860: inst = 32'h00000000;
32'd864: inst = 32'h080000d6;
32'd868: inst = 32'h00000000;
32'd872: inst = 32'h00000000;
32'd876: inst = 32'h20080380;
32'd880: inst = 32'h01000008;
32'd884: inst = 32'h00000000;
32'd888: inst = 32'h080000de;
32'd892: inst = 32'h00000000;
32'd896: inst = 32'h00000000;
32'd900: inst = 32'h20080398;
32'd904: inst = 32'h0100f809;
32'd908: inst = 32'h00000000;
32'd912: inst = 32'h080000e4;
32'd916: inst = 32'h00000000;
32'd920: inst = 32'h200f0390;
32'd924: inst = 32'h17effffe;
32'd928: inst = 32'h00000000;
32'd932: inst = 32'h00000000;
32'd936: inst = 32'h20080000;
32'd940: inst = 32'h2009ffff;
32'd944: inst = 32'h0109502a;
32'd948: inst = 32'h0128582b;
32'd952: inst = 32'h1540ffff;
32'd956: inst = 32'h00000000;
32'd960: inst = 32'h1560fffd;
32'd964: inst = 32'h00000000;
32'd968: inst = 32'h00000000;
32'd972: inst = 32'h20080001;
32'd976: inst = 32'h2009ffff;
32'd980: inst = 32'h01095024;
32'd984: inst = 32'h01095825;
32'd988: inst = 32'h01096026;
32'd992: inst = 32'h01096827;
32'd996: inst = 32'h200f0001;
32'd1000: inst = 32'h154ffffe;
32'd1004: inst = 32'h00000000;
32'd1008: inst = 32'h200fffff;
32'd1012: inst = 32'h156ffffb;
32'd1016: inst = 32'h00000000;
32'd1020: inst = 32'h200ffffe;
32'd1024: inst = 32'h158ffff8;
32'd1028: inst = 32'h00000000;
32'd1032: inst = 32'h200f0000;
32'd1036: inst = 32'h15affff5;
32'd1040: inst = 32'h00000000;
32'd1044: inst = 32'h00000000;
32'd1048: inst = 32'h20080001;
32'd1052: inst = 32'h2009ffff;
32'd1056: inst = 32'h01095022;
32'd1060: inst = 32'h01095823;
32'd1064: inst = 32'h200f0002;
32'd1068: inst = 32'h154ffffe;
32'd1072: inst = 32'h00000000;
32'd1076: inst = 32'h156ffffc;
32'd1080: inst = 32'h00000000;
32'd1084: inst = 32'h00000000;
32'd1088: inst = 32'h20080001;
32'd1092: inst = 32'h2009ffff;
32'd1096: inst = 32'h01095020;
32'd1100: inst = 32'h01095821;
32'd1104: inst = 32'h1540ffff;
32'd1108: inst = 32'h00000000;
32'd1112: inst = 32'h1560fffd;
32'd1116: inst = 32'h00000000;
32'd1120: inst = 32'h00000000;
32'd1124: inst = 32'h20080003;
32'd1128: inst = 32'h2009fffe;
32'd1132: inst = 32'h0109001b;
32'd1136: inst = 32'h00000000;
32'd1140: inst = 32'h00005010;
32'd1144: inst = 32'h200f0003;
32'd1148: inst = 32'h154ffffc;
32'd1152: inst = 32'h00000000;
32'd1156: inst = 32'h00000000;
32'd1160: inst = 32'h00005012;
32'd1164: inst = 32'h1540fffd;
32'd1168: inst = 32'h00000000;
32'd1172: inst = 32'h00000000;
32'd1176: inst = 32'h20080003;
32'd1180: inst = 32'h2009fffe;
32'd1184: inst = 32'h0109001a;
32'd1188: inst = 32'h00000000;
32'd1192: inst = 32'h00005010;
32'd1196: inst = 32'h200f0001;
32'd1200: inst = 32'h154ffffc;
32'd1204: inst = 32'h00000000;
32'd1208: inst = 32'h00000000;
32'd1212: inst = 32'h00005012;
32'd1216: inst = 32'h200fffff;
32'd1220: inst = 32'h154ffffc;
32'd1224: inst = 32'h00000000;
32'd1228: inst = 32'h00000000;
32'd1232: inst = 32'h2008ffff;
32'd1236: inst = 32'h2009ffff;
32'd1240: inst = 32'h01090019;
32'd1244: inst = 32'h00005010;
32'd1248: inst = 32'h214a0002;
32'd1252: inst = 32'h1540fffd;
32'd1256: inst = 32'h00000000;
32'd1260: inst = 32'h00000000;
32'd1264: inst = 32'h00005012;
32'd1268: inst = 32'h200f0001;
32'd1272: inst = 32'h154ffffc;
32'd1276: inst = 32'h00000000;
32'd1280: inst = 32'h00000000;
32'd1284: inst = 32'h2008ffff;
32'd1288: inst = 32'h2009ffff;
32'd1292: inst = 32'h01090018;
32'd1296: inst = 32'h00005010;
32'd1300: inst = 32'h1540fffe;
32'd1304: inst = 32'h00000000;
32'd1308: inst = 32'h00000000;
32'd1312: inst = 32'h00005012;
32'd1316: inst = 32'h200f0001;
32'd1320: inst = 32'h154ffffc;
32'd1324: inst = 32'h00000000;
32'd1328: inst = 32'h00000000;
32'd1332: inst = 32'h20080001;
32'd1336: inst = 32'h01000013;
32'd1340: inst = 32'h00004812;
32'd1344: inst = 32'h200f0001;
32'd1348: inst = 32'h152ffffe;
32'd1352: inst = 32'h00000000;
32'd1356: inst = 32'h00000000;
32'd1360: inst = 32'h20080001;
32'd1364: inst = 32'h01000011;
32'd1368: inst = 32'h00004810;
32'd1372: inst = 32'h200f0001;
32'd1376: inst = 32'h152ffffe;
32'd1380: inst = 32'h00000000;
32'd1384: inst = 32'h00000000;
32'd1388: inst = 32'h20080001;
32'd1392: inst = 32'h00084840;
32'd1396: inst = 32'h200f0002;
32'd1400: inst = 32'h152ffffe;
32'd1404: inst = 32'h00000000;
32'd1408: inst = 32'h00000000;
32'd1412: inst = 32'h20080002;
32'd1416: inst = 32'h00084842;
32'd1420: inst = 32'h200f0001;
32'd1424: inst = 32'h152ffffe;
32'd1428: inst = 32'h00000000;
32'd1432: inst = 32'h00000000;
32'd1436: inst = 32'h20080000;
32'd1440: inst = 32'h20090001;
32'd1444: inst = 32'h01094022;
32'd1448: inst = 32'h00085043;
32'd1452: inst = 32'h1548ffff;
32'd1456: inst = 32'h00000000;
32'd1460: inst = 32'h00000000;
32'd1464: inst = 32'h20080001;
32'd1468: inst = 32'h20090003;
32'd1472: inst = 32'h01285004;
32'd1476: inst = 32'h200f0008;
32'd1480: inst = 32'h154ffffe;
32'd1484: inst = 32'h00000000;
32'd1488: inst = 32'h00000000;
32'd1492: inst = 32'h20080000;
32'd1496: inst = 32'h20090001;
32'd1500: inst = 32'h01094022;
32'd1504: inst = 32'h200a0003;
32'd1508: inst = 32'h01485007;
32'd1512: inst = 32'h1548ffff;
32'd1516: inst = 32'h00000000;
		
			default: 	inst = 32'hxxxxxxxx;
		endcase
	end

endmodule
